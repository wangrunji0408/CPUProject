library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Base.all;

-- 取指模块
entity IF_ is
	port (
		rst, clk: in std_logic
	) ;
end IF_;

architecture arch of IF_ is	
begin

end arch ; -- arch
