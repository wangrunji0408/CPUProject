library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Base.all;

-- 寄存器堆
entity Register is
	port (
		clk, rst: in std_logic;
		write: in RegPort;
		read1, read2: inout RegPort -- only .data is out
	) ;
end Register;

architecture arch of Register is	
begin
	-- 1. $0=0
	-- 2. 读使能无效时，输出0
	-- 3. 时钟上升沿时，若写使能生效，将数据写入
end arch ; -- arch
